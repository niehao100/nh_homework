`timescale 1ns/1ps
module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];
localparam ROM_SIZE = 32;
always@(*)
    case(addr)	//Address Must Be Word Aligned.
32'b00000000000000000000000000000000: data <= 32'b00111100000101010100000000000000;// lui $s5,16384
32'b00000000000000000000000000000100: data <= 32'b00100000000010010000000000000000;// addi $t1,$zero, 0
32'b00000000000000000000000000001000: data <= 32'b10101110101010010000000000001000;// sw $t1,8($s5)
32'b00000000000000000000000000001100: data <= 32'b00100000000001010000000100000000;// addi $a1,$zero, 256
32'b00000000000000000000000000010000: data <= 32'b00100000000010010000000000000100;// addi $t1,$zero, 4
32'b00000000000000000000000000010100: data <= 32'b10101110101010010000000000100000;// sw $t1,32($s5)
// Loop1:
32'b00000000000000000000000000011000: data <= 32'b10001110101000100000000000011100;// lw $v0,28($s5)
32'b00000000000000000000000000011100: data <= 32'b00010000010000001111111111111110;// beq $v0,$zero, Loop1
32'b00000000000000000000000000100000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000000100100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000000101000: data <= 32'b00100000000010010000000000000000;// addi $t1,$zero, 0
32'b00000000000000000000000000101100: data <= 32'b10101110101010010000000000100000;// sw $t1,32($s5)
32'b00000000000000000000000000110000: data <= 32'b00000000000000101000100000100000;// add $s1,$zero, $v0
32'b00000000000000000000000000110100: data <= 32'b10101110101000100000000000001100;// sw $v0,12($s5)
32'b00000000000000000000000000111000: data <= 32'b00100000000010110000000000000001;// addi $t3,$zero, 1
32'b00000000000000000000000000111100: data <= 32'b00100000000010100000000110010000;// addi $t2,$zero, 400
// L2:
32'b00000000000000000000000001000000: data <= 32'b00000001010010110101000000100010;// sub $t2,$t2, $t3
32'b00000000000000000000000001000100: data <= 32'b00010101010000001111111111111110;// bne $t2,$zero, L2
32'b00000000000000000000000001001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000001001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000001010000: data <= 32'b00100000000010010000000000000100;// addi $t1,$zero, 4
32'b00000000000000000000000001010100: data <= 32'b10101110101010010000000000100000;// sw $t1,32($s5)
// Loop2:
32'b00000000000000000000000001011000: data <= 32'b10001110101000110000000000011100;// lw $v1,28($s5)
32'b00000000000000000000000001011100: data <= 32'b00010000011000001111111111111110;// beq $v1,$zero, Loop2
32'b00000000000000000000000001100000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000001100100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000001101000: data <= 32'b00100000000010010000000000000000;// addi $t1,$zero, 0
32'b00000000000000000000000001101100: data <= 32'b10101110101010010000000000100000;// sw $t1,32($s5)
32'b00000000000000000000000001110000: data <= 32'b00000000000000111001000000100000;// add $s2,$zero, $v1
32'b00000000000000000000000001110100: data <= 32'b10101110101000110000000000001100;// sw $v1,12($s5)
32'b00000000000000000000000001111000: data <= 32'b00100000000010100010011100010000;// addi $t2,$zero, 10000
// L4:
32'b00000000000000000000000001111100: data <= 32'b00000001010010110101000000100010;// sub $t2,$t2, $t3
32'b00000000000000000000000010000000: data <= 32'b00010101010000001111111111111110;// bne $t2,$zero, L4
32'b00000000000000000000000010000100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000010001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000010001100: data <= 32'b00000000000000100001001000000000;// sll $v0,$v0, 8
32'b00000000000000000000000010010000: data <= 32'b00000000010000110001100000100000;// add $v1,$v0, $v1
32'b00000000000000000000000010010100: data <= 32'b00010010001100100000000000001110;// beq $s1,$s2, output
32'b00000000000000000000000010011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000010011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// judge:
32'b00000000000000000000000010100000: data <= 32'b00000010010100010100100000100010;// sub $t1,$s2, $s1
32'b00000000000000000000000010100100: data <= 32'b00011001001000000000000000000101;// blez $t1,loop3
32'b00000000000000000000000010101000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000010101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// bigger:
32'b00000000000000000000000010110000: data <= 32'b00100010010010010000000000000000;// addi $t1,$s2, 0
32'b00000000000000000000000010110100: data <= 32'b00100010001100100000000000000000;// addi $s2,$s1, 0
32'b00000000000000000000000010111000: data <= 32'b00100001001100010000000000000000;// addi $s1,$t1, 0
// loop3:
32'b00000000000000000000000010111100: data <= 32'b00000010001100101001100000100010;// sub $s3,$s1, $s2
32'b00000000000000000000000011000000: data <= 32'b00100010011100010000000000000000;// addi $s1,$s3, 0
32'b00000000000000000000000011000100: data <= 32'b00010110001100101111111111110110;// bne $s1,$s2, judge
32'b00000000000000000000000011001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000011001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// output:
32'b00000000000000000000000011010000: data <= 32'b00100000000010010000000000000001;// addi $t1,$zero, 1
32'b00000000000000000000000011010100: data <= 32'b10101110101100010000000000011000;// sw $s1,24($s5)
32'b00000000000000000000000011011000: data <= 32'b10101110101100010000000000001100;// sw $s1,12($s5)
32'b00000000000000000000000011011100: data <= 32'b00000000000010010101000000100010;// sub  $t2,$zero, $t1
32'b00000000000000000000000011100000: data <= 32'b10101110101010100000000000000100;// sw $t2,4($s5)
32'b00000000000000000000000011100100: data <= 32'b00100000000011000000000001100100;// addi $t4,$zero, 100 
32'b00000000000000000000000011101000: data <= 32'b00000001010011000101100000100010;// sub $t3,$t2, $t4 
32'b00000000000000000000000011101100: data <= 32'b10101110101010110000000000000000;// sw $t3,0($s5)
32'b00000000000000000000000011110000: data <= 32'b00100000000010100000000000000011;// addi $t2,$zero, 3
32'b00000000000000000000000011110100: data <= 32'b00100000000000100000000000000001;// addi $v0,$zero, 1
32'b00000000000000000000000011111000: data <= 32'b10101110101010100000000000001000;// sw $t2,8($s5)
32'b00000000000000000000000011111100: data <= 32'b00000000000011000010000000100000;// add $a0,$zero, $t4
// LOOP4:
32'b00000000000000000000000100000000: data <= 32'b00100000000100100000000000000000;// addi $s2,$zero, 0 
32'b00000000000000000000000100000100: data <= 32'b00001000000000000000000001000000;// j LOOP4
32'b00000000000000000000000100001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b00000000000000000000000100001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// DECODE:
32'b10000000000000000000000100010000: data <= 32'b00100000000010110000000010000000;// addi $t3,$zero, 128
32'b10000000000000000000000100010100: data <= 32'b00100000011011010000000000000000;// addi $t5,$v1, 0
// SHIFTL:
32'b10000000000000000000000100011000: data <= 32'b00010001011000100000000000000111;// beq $t3,$v0, SHIFTR
32'b10000000000000000000000100011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000100100000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000100100100: data <= 32'b00000000000011010110100100000000;// sll $t5,$t5, 4
32'b10000000000000000000000100101000: data <= 32'b00000000000010110101100001000010;// srl $t3,$t3, 1
32'b10000000000000000000000100101100: data <= 32'b00001000000000000000000001000110;// j SHIFTL
32'b10000000000000000000000100110000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000100110100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// SHIFTR:
32'b10000000000000000000000100111000: data <= 32'b00000000000011010110111100000010;// srl $t5,$t5, 28
32'b10000000000000000000000100111100: data <= 32'b00000000000010110101101000000000;// sll $t3,$t3, 8
32'b10000000000000000000000101000000: data <= 32'b00100000000011100000000000000000;// addi $t6,$zero, 0
32'b10000000000000000000000101000100: data <= 32'b00010001110011010000000000111110;// beq $t6,$t5, ZERO
32'b10000000000000000000000101001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101010000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000101010100: data <= 32'b00010001110011010000000000111100;// beq $t6,$t5, ONE
32'b10000000000000000000000101011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101100000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000101100100: data <= 32'b00010001110011010000000000111010;// beq $t6,$t5, TWO
32'b10000000000000000000000101101000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101110000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000101110100: data <= 32'b00010001110011010000000000111000;// beq $t6,$t5, THREE
32'b10000000000000000000000101111000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000101111100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110000000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000110000100: data <= 32'b00010001110011010000000000110110;// beq $t6,$t5, FOUR
32'b10000000000000000000000110001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110010000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000110010100: data <= 32'b00010001110011010000000000110100;// beq $t6,$t5, FIVE
32'b10000000000000000000000110011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110100000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000110100100: data <= 32'b00010001110011010000000000110010;// beq $t6,$t5, SIX
32'b10000000000000000000000110101000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110110000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000110110100: data <= 32'b00010001110011010000000000110000;// beq $t6,$t5, SEVEN
32'b10000000000000000000000110111000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000110111100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111000000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000111000100: data <= 32'b00010001110011010000000000101110;// beq $t6,$t5, EIGHT
32'b10000000000000000000000111001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111010000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000111010100: data <= 32'b00010001110011010000000000101100;// beq $t6,$t5, NIGHT
32'b10000000000000000000000111011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111100000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000111100100: data <= 32'b00010001110011010000000000101010;// beq $t6,$t5, A
32'b10000000000000000000000111101000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111110000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000000111110100: data <= 32'b00010001110011010000000000101000;// beq $t6,$t5, B
32'b10000000000000000000000111111000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000111111100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000000000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000001000000100: data <= 32'b00010001110011010000000000100110;// beq $t6,$t5, C
32'b10000000000000000000001000001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000010000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000001000010100: data <= 32'b00010001110011010000000000100100;// beq $t6,$t5, D
32'b10000000000000000000001000011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000011100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000100000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000001000100100: data <= 32'b00010001110011010000000000100010;// beq $t6,$t5, E
32'b10000000000000000000001000101000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000110000: data <= 32'b00100001110011100000000000000001;// addi $t6,$t6, 1
32'b10000000000000000000001000110100: data <= 32'b00010001110011010000000000100000;// beq $t6,$t5, F
32'b10000000000000000000001000111000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001000111100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// ZERO:
32'b10000000000000000000001001000000: data <= 32'b00100000000011010000000001000000;// addi $t5,$zero, 64
32'b10000000000000000000001001000100: data <= 32'b00001000000000000000000010110000;// j DE
// ONE:
32'b10000000000000000000001001001000: data <= 32'b00100000000011010000000001111001;// addi $t5,$zero, 121
32'b10000000000000000000001001001100: data <= 32'b00001000000000000000000010110000;// j DE
// TWO:
32'b10000000000000000000001001010000: data <= 32'b00100000000011010000000000100100;// addi $t5,$zero, 36
32'b10000000000000000000001001010100: data <= 32'b00001000000000000000000010110000;// j DE
// THREE:
32'b10000000000000000000001001011000: data <= 32'b00100000000011010000000000110000;// addi $t5,$zero, 48
32'b10000000000000000000001001011100: data <= 32'b00001000000000000000000010110000;// j DE
// FOUR:
32'b10000000000000000000001001100000: data <= 32'b00100000000011010000000000011001;// addi $t5,$zero, 25
32'b10000000000000000000001001100100: data <= 32'b00001000000000000000000010110000;// j DE
// FIVE:
32'b10000000000000000000001001101000: data <= 32'b00100000000011010000000000010010;// addi $t5,$zero, 18
32'b10000000000000000000001001101100: data <= 32'b00001000000000000000000010110000;// j DE
// SIX:
32'b10000000000000000000001001110000: data <= 32'b00100000000011010000000000000010;// addi $t5,$zero, 2
32'b10000000000000000000001001110100: data <= 32'b00001000000000000000000010110000;// j DE
// SEVEN:
32'b10000000000000000000001001111000: data <= 32'b00100000000011010000000001111000;// addi $t5,$zero, 120
32'b10000000000000000000001001111100: data <= 32'b00001000000000000000000010110000;// j DE
// EIGHT:
32'b10000000000000000000001010000000: data <= 32'b00100000000011010000000000000000;// addi $t5,$zero, 0
32'b10000000000000000000001010000100: data <= 32'b00001000000000000000000010110000;// j DE
// NIGHT:
32'b10000000000000000000001010001000: data <= 32'b00100000000011010000000000010000;// addi $t5,$zero, 16
32'b10000000000000000000001010001100: data <= 32'b00001000000000000000000010110000;// j DE
// A:
32'b10000000000000000000001010010000: data <= 32'b00100000000011010000000000001000;// addi $t5,$zero, 8
32'b10000000000000000000001010010100: data <= 32'b00001000000000000000000010110000;// j DE
// B:
32'b10000000000000000000001010011000: data <= 32'b00100000000011010000000000000011;// addi $t5,$zero, 3
32'b10000000000000000000001010011100: data <= 32'b00001000000000000000000010110000;// j DE
// C:
32'b10000000000000000000001010100000: data <= 32'b00100000000011010000000001000110;// addi $t5,$zero, 70
32'b10000000000000000000001010100100: data <= 32'b00001000000000000000000010110000;// j DE
// D:
32'b10000000000000000000001010101000: data <= 32'b00100000000011010000000000100001;// addi $t5,$zero, 33
32'b10000000000000000000001010101100: data <= 32'b00001000000000000000000010110000;// j DE
// E:
32'b10000000000000000000001010110000: data <= 32'b00100000000011010000000000000110;// addi $t5,$zero, 6
32'b10000000000000000000001010110100: data <= 32'b00001000000000000000000010110000;// j DE
// F:
32'b10000000000000000000001010111000: data <= 32'b00100000000011010000000000001110;// addi $t5,$zero, 14
32'b10000000000000000000001010111100: data <= 32'b00001000000000000000000010110000;// j DE
// DE:
32'b10000000000000000000001011000000: data <= 32'b00000001011011010110100000100000;// add $t5,$t3, $t5
32'b10000000000000000000001011000100: data <= 32'b10101110101011010000000000010100;// sw $t5,20($s5)
32'b10000000000000000000001011001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011010000: data <= 32'b00000000000000100001000001000000;// sll $v0,$v0, 1
32'b10000000000000000000001011010100: data <= 32'b00100000000010110000000000010000;// addi $t3,$zero, 16
32'b10000000000000000000001011011000: data <= 32'b00100000000010010000000000000011;// addi $t1,$zero, 3
32'b10000000000000000000001011011100: data <= 32'b10101110101010010000000000001000;// sw $t1,8($s5)
32'b10000000000000000000001011100000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011100100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011101000: data <= 32'b00010100010010110000000000000101;// bne $v0,$t3, JUMP
32'b10000000000000000000001011101100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011110000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011110100: data <= 32'b00100000000000100000000000000001;// addi $v0,$zero, 1
32'b10000000000000000000001011111000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001011111100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
// JUMP:
32'b10000000000000000000001100000000: data <= 32'b00000000101000000000000000001000;// jr $a1
32'b10000000000000000000001100000100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001100001000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000001100001100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000000000100: data <= 32'b00100000000010010000000000000001;// addi $t1,$zero, 0
32'b10000000000000000000000000001000: data <= 32'b10101110101010010000000000001000;// sw $t1,8($s5)
32'b10000000000000000000000000001100: data <= 32'b00001100000000000000000001000100;// jal DECODE
32'b10000000000000000000000000010000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000000010100: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0
32'b10000000000000000000000000011000: data <= 32'b00000000000000000000000000000000;// sll $zero,$zero, 0

        default:	data <= 32'h0000_0008;
endcase
endmodule