`timescale 1ns/1ps
module ROM (addr,data,enable);
input [31:0] addr;
input enable;
output [31:0] data;
reg [31:0] tempdata;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];
assign data=enable? tempdata : 32'b0;
always@(*)
    case(addr)	//Address Must Be Word Aligned.
32'b00000000000000000000000000000000: tempdata <= 32'b00111100000101010100000000000000;// lui $s5,16384
32'b00000000000000000000000000000100: tempdata <= 32'b00100000000010010000000000000000;// addi $t1,$zero, 0
32'b00000000000000000000000000001000: tempdata <= 32'b10101110101010010000000000001000;// sw $t1,8($s5)
// L1:
32'b00000000000000000000000000001100: tempdata <= 32'b10001110101000100000000000011100;// lw $v0,28($s5)
32'b00000000000000000000000000010000: tempdata <= 32'b00010000010010011111111111111110;// beq $v0,$t1, L1
32'b00000000000000000000000000010100: tempdata <= 32'b00000000000000101000100000100000;// add $s1,$zero, $v0
32'b00000000000000000000000000011000: tempdata <= 32'b10101110101100010000000000011000;// sw $s1,24($s5)
32'b00000000000000000000000000011100: tempdata <= 32'b00100000000010100010011100010000;// addi $t2,$zero, 10000
32'b00000000000000000000000000100000: tempdata <= 32'b00100000000010110000000000000001;// addi $t3,$zero, 1
// LOOP:
32'b00000000000000000000000000100100: tempdata <= 32'b00000001010010110101000000100010;// sub $t2,$t2, $t3
32'b00000000000000000000000000101000: tempdata <= 32'b00010101010010011111111111111110;// bne $t2,$t1, LOOP
32'b00000000000000000000000000101100: tempdata <= 32'b00001000000000000000000000000011;// j L1

        default:	tempdata <= 32'h0000_0008;
endcase
endmodule