`timescale 1ns/1ps
//modefied by Neil

module Peripheral (reset,clk,rd,wr,addr,wdata,rdata,led,switch,digi,irqout);

input reset,clk;
input rd,wr;
input [31:0] addr;
input [31:0] wdata;
input [7:0] switch;

output  irqout;
output [7:0] led;
output [11:0] digi;
output [31:0] rdata;

reg [2:0] TCON;
reg [7:0] led;
reg [11:0] digi;
reg [31:0] TH,TL;
reg [31:0] rdata;

initial begin
    TCON=3'b000;
	digi=11'b0;
	led=8'b0;
end
assign irqout = TCON[2];

	


always@(*) begin
	if(rd) begin
		case(addr)
			32'h40000000: rdata<=TH;			
			32'h40000004: rdata<=TL;			
			32'h40000008: rdata<={29'b0,TCON};				
			32'h4000000C: rdata<={24'b0,led};			
			32'h40000010: rdata<={24'b0,switch};
			32'h40000014: rdata<={20'b0,digi};
			default: rdata<=32'b0;
		endcase
	end
	else
		rdata<=32'b0;
end


always@(negedge reset or posedge clk) begin
	if(~reset) begin
		TH<=32'b0;
		TL<=32'b0;
		TCON<=3'b0;
		led<=8'b0;
		digi<=12'b0;	
	end
	else begin
		if(TCON[0]) begin	//timer is enabled
			if(TL==32'hffffffff) begin
				TL<=TH;
				if(TCON[1]) TCON<=3'b101;		//irq is enabled
			end
            else begin
                TL<=TL + 1;
                TCON[2]<=1'b0;
            end
		end
		
		if(wr) begin
			case(addr)
				32'h40000000: TH<=wdata;
				32'h40000004: TL<=wdata;
				32'h40000008: TCON<=wdata[2:0];		
				32'h4000000C: led<=wdata[7:0];			
				32'h40000014: digi<=wdata[11:0];
				default: ;
			endcase
		end
	end
end
endmodule

